`timescale 1 ns/10 ps  // time-unit = 1 ns, precision = 10 ps

// dummy implementation, please replace with your own
module sequential_circuits ( 
    input clk,    // Clocks are used in sequential circuits
    input d,
    output q );//



    assign q = d;

endmodule